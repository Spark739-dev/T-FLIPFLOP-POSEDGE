library verilog;
use verilog.vl_types.all;
entity tfliflop_vlg_vec_tst is
end tfliflop_vlg_vec_tst;
